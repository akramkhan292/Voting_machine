/home/nilet/akram/voting_machine/counter_design_database_45nm/lef/gsclib045_tech.lef